initial begin
  ascend = '{0,1,2,3};
  $display("%p", ascend);
end
